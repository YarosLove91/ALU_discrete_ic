// Модель микросхемы 74882 - микросхема ускоренного переноса (CLA) на 32 бита.
// Для работы требуется 8 битный сумматор или АЛУ

module cla32_n74882 (
    input [7:0] nP,      // Пропускные сигналы
    input [7:0] nG,      // Генерирующие сигналы
    input Cin,           // Входной перенос
    output Cn_8, Cn_16, Cn_24, Cn_32    // Выходные переносы
);
    // Используется компактная форма записи
    // Активный уровень - 0
    assign Cn_8 = ~((nG[1] & nP[1]) | 
                      (&(nG[1:0]) & nP[0])| 
                      (&(nG[1:0]) & ~Cin));
    
    assign Cn_16 = ~ ((nG[3] & nP[3]) | 
                       (&(nG[3:2]) & nP[2]) |
                       (&(nG[3:1]) & nP[1]) |
                       (&(nG[3:0]) & nP[0]) |
                       (&(nG[3:0]) & ~Cin));

    assign Cn_24 = ~((nG[5] & nP[5]) |
                      (&(nG[5:4]) & nP[4]) |
                      (&(nG[5:3]) & nP[3]) |
                      (&(nG[5:2]) & nP[2]) |
                      (&(nG[5:1]) & nP[1]) |
                      (&(nG[5:0]) & nP[0]) |
                      (&(nG[5:0]) & ~Cin));

    assign Cn_32 = ~((nG[7] & nP[7]) |
                      (&(nG[7:6]) & nP[6]) |
                      (&(nG[7:5]) & nP[5]) |
                      (&(nG[7:4]) & nP[4]) |
                      (&(nG[7:3]) & nP[3]) |
                      (&(nG[7:2]) & nP[2]) |
                      (&(nG[7:1]) & nP[1]) |
                      (&(nG[7:0]) & nP[0]) |
                      (&(nG[7:0]) & ~Cin));

endmodule 